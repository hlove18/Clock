include 
begin
end
fork

addc
add 
ajmp
sjmp
anl

